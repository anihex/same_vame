module main

fn main() {
	println('Hello World !')
}
